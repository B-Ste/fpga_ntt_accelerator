`timescale 1ns/1ps

module modular_multiplier_tb ();

    reg clk = 0;
    reg [29:0]a;
    reg [29:0]b;
    wire [29:0]c;

    modular_multiplier #12 mult (clk, a, b, c);

    always #50 clk = ~clk;

    initial
    begin
        a <= 100;
        b <= 1000;
        #100;
        a <= 12345;
        b <= 12345;
        #100;
        a <= 9582;
        b <= 6847912;
        #100;
        a <= 1063321600;
        b <= 1063321600;
        #100;
        a <= 1063452672;
        b <= 1063452672;
        #100;
        a <= 1064697856;
        b <= 1064697856;
        #100;
        a <= 1065484288;
        b <= 1065484288;
        #100;
        a <= 1065811968;
        b <= 1065811968;
        #100; 
        a <= 1068236800;
        b <= 1068236800;
        #100;
        a <= 1068433408;
        b <= 1068433408;
        #100;
        a <= 1068564480;
        b <= 1068564480;
        #100;
        a <= 1069219840;
        b <= 1069219840;
        #100;
        a <= 1070727168;
        b <= 1070727168;
        #100;
        a <= 1071513600;
        b <= 1071513600;
        #100;
        a <= 1072496640;
        b <= 1072496640;
        #100;
        a <= 1073479680;
        b <= 1073479680;
        #1000;
    end
    
endmodule
